
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity stock is
    generic (
        NUM_PRODUCTOS : positive := 9;
        PROD_BITS     : positive := 4   -- permite codificar hasta 9 productos
    );
    port(
        clk             : in  std_logic;
        estado          : in  unsigned(2 downto 0);
        productos       : in  std_logic_vector(NUM_PRODUCTOS-1 downto 0);
        error_pago      : in  std_logic;
        RESET_STOCK     : in  std_logic;
        Boton_Confirmar : in  std_logic;
        
        productoOk     : out std_logic;
        errorProducto  : out std_logic;
        producto_id    : out unsigned(PROD_BITS-1 downto 0);  --prod. determinista 
        STOCK_producto_i   : out std_logic_vector(NUM_PRODUCTOS-1 downto 0)
    );
end stock;

architecture Behavioral of stock is

    -- memoria de stock (9 productos)
    type stock_array_t is array (0 to NUM_PRODUCTOS-1) of unsigned(3 downto 0);

    -- Valores "de fabrica" para poder restaurar con RESET_STOCK
    constant STOCK_INIT : stock_array_t := (
        to_unsigned(5,4),  -- producto 0
        to_unsigned(3,4),  -- producto 1
        to_unsigned(7,4),  -- producto 2
        to_unsigned(3,4),  -- producto 3
        to_unsigned(4,4),  -- producto 4
        to_unsigned(6,4),  -- producto 5
        to_unsigned(3,4),  -- producto 6
        to_unsigned(8,4),  -- producto 7
        to_unsigned(9,4)   -- producto 8
    );

    constant ESTADO_0 : unsigned(2 downto 0) := (others => '0');             

    signal stock_mem        : stock_array_t := STOCK_INIT;                      -- INICIALIZACION A VALORES POR DEFECTO stock

    signal productoOk_reg     : std_logic := '0';
    signal errorProducto_reg  : std_logic := '0';

    signal idx               : integer range 0 to NUM_PRODUCTOS-1 := 0;
    signal seleccion_valida  : std_logic := '0';  -- exactamente un bit a '1'
    
    -- Combinacional: validar one-hot y extraer indice
    signal prod_u        : unsigned(NUM_PRODUCTOS-1 downto 0);
    signal onehot_valid  : std_logic;
    signal sel_idx       : unsigned(PROD_BITS-1 downto 0);

    signal producto_id_reg   : unsigned(PROD_BITS-1 downto 0);  --prod. determinista 
    signal estado_prev       : unsigned(2 downto 0) := (others => '0');

    signal stock_bar_reg : std_logic_vector(NUM_PRODUCTOS-1 downto 0) := (others => '0');

begin

    prod_u <= unsigned(productos);

    -- onehot_valid = (productos != 0) AND ((productos AND (productos-1)) = 0)
    onehot_valid <= '1' when (prod_u /= 0) and ((prod_u and (prod_u - 1)) = 0) else '0';

    -- Decodificar indice (combinacional, simple)
    process(prod_u)
        variable tmp : unsigned(PROD_BITS-1 downto 0);
    begin
        tmp := (others => '0');
        for i in 0 to NUM_PRODUCTOS-1 loop
            if prod_u(i) = '1' then
                tmp := to_unsigned(i, PROD_BITS);
            end if;
        end loop;
        sel_idx <= tmp;
    end process;
----------------------------------------------------------

-- Ejemplos (NUM_PRODUCTOS=9): 0->000000000, 1->100000000, 2->110000000, 3->111000000, 7->111111100
process(onehot_valid, sel_idx)
    variable nn : integer;
begin
    stock_bar_reg <= (others => '0');
    nn := 0;

    if onehot_valid = '1' then
        nn := to_integer(stock_mem(to_integer(sel_idx)));

        -- Saturar por si el stock fuese mayor que NUM_PRODUCTOS
        if nn > NUM_PRODUCTOS then
            nn := NUM_PRODUCTOS;
        elsif nn < 0 then
            nn := 0;
        end if;

        -- Bucle de rango CONSTANTE (sintetizable)
        for k in 0 to NUM_PRODUCTOS-1 loop
            if k < nn then
                stock_bar_reg(NUM_PRODUCTOS-1-k) <= '1';  -- barra desde MSB
            end if;
        end loop;
    end if;
end process;





-------------------------------------------------------
    -- Secuencial
    process(clk)
    begin

      if rising_edge(clk) then
    
        -- Pulsos por defecto (1 ciclo)
        productoOk_reg    <= '0';
        errorProducto_reg <= '0';
    
        -- Detectar re-entrada en estado 0 para limpiar lo mostrado
        if (estado_prev /= ESTADO_0) and (estado = ESTADO_0) then
          producto_id_reg <= to_unsigned(0, PROD_BITS);
        end if;
        estado_prev <= estado;
    
        -- Reset del stock a valores de fabrica                         -- HE CAMBIADO EL RESET A 0
        if RESET_STOCK = '0' then
          stock_mem       <= STOCK_INIT;
          producto_id_reg <= to_unsigned(0, PROD_BITS);
    
        else
          -- Solo trabajamos en estado 0
          if estado = ESTADO_0 then
    
            -- Si hay error de pago: bloqueo total (no comprar, no tocar stock)
            if error_pago = '1' then
              -- si quieres que no se muestre ningun producto cuando hay error de pago:
              producto_id_reg <= to_unsigned(0, PROD_BITS);
    
            else
              -- Solo actuamos si confirman (idealmente esto es un pulso)
              if Boton_Confirmar = '1' then
    
                -- Seleccion invalida (ninguno o varios) => errorProducto
                if onehot_valid = '0' then
                  errorProducto_reg <= '1';
                else
                  -- Seleccion valida: mirar stock
                  if stock_mem(to_integer(sel_idx)) > 0 then
                    stock_mem(to_integer(sel_idx)) <= stock_mem(to_integer(sel_idx)) - 1;
                    productoOk_reg  <= '1';
                    producto_id_reg <= sel_idx;
                  else
                    errorProducto_reg <= '1';
                  end if;
                end if;
              end if;
            end if;
          end if;
        end if;

  end if;
end process;

    productoOk    <= productoOk_reg;
    errorProducto <= errorProducto_reg;
    producto_id   <= producto_id_reg;
    
    
    -- Barra de bits de stock por producto seleccionado
    STOCK_producto_i <= stock_bar_reg;

end Behavioral;





library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity SINCRONIZADOR is
    generic(
        NUM_MONEDAS: positive:= 4;
        NUM_PRODUCTOS: positive:= 9
    );
    
    port(
        CLK: in std_logic;

        AS_PRODUCTOS: in std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
        AS_MONEDAS: in std_logic_vector (NUM_MONEDAS - 1 downto 0); 
        AS_CONFI : in std_logic;
    
        S_PRODUCTOS: out std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
        S_MONEDAS: out std_logic_vector (NUM_MONEDAS - 1 downto 0);
        S_CONFI : out std_logic

    );   
    
         
end SINCRONIZADOR;

architecture Behavioral of SINCRONIZADOR is

    signal REG1_PRODUCTOS: std_logic_vector (NUM_PRODUCTOS - 1 downto 0);    
    signal REG1_MONEDAS: std_logic_vector(NUM_MONEDAS - 1 downto 0);
    signal REG1_CONFI: std_logic;

    signal REG2_PRODUCTOS: std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
    signal REG2_MONEDAS: std_logic_vector(NUM_MONEDAS - 1 downto 0);
    signal REG2_CONFI: std_logic;  

begin

    REGISTRO_1: process(CLK)
    begin
        if rising_edge(CLK) then
            REG1_PRODUCTOS<= AS_PRODUCTOS;
            REG1_MONEDAS<= AS_MONEDAS;
            REG1_CONFI <= AS_CONFI;
            
        end if;
    end process;
    
    REGISTRO_2:process(CLK)
    begin
        if rising_edge(CLK) then
            REG2_PRODUCTOS<= REG1_PRODUCTOS;        
            REG2_MONEDAS<= REG1_MONEDAS;
            REG2_CONFI <= REG1_CONFI;
        end if;
    end process;

    S_MONEDAS <= REG2_MONEDAS;
    S_PRODUCTOS<= REG2_PRODUCTOS;
    S_CONFI <= REG2_CONFI;
    
end Behavioral;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TOP is
generic (
        Monedas       : POSITIVE := 4;   -- genérico con valor por defecto 4
        NUM_PRODUCTOS : POSITIVE := 9;   -- genérico con valor por defecto 9
        NUM_DIGITS    : positive := 8;
        NUM_SEGS      : positive := 8;   -- antes 7, ahora 8 (anodos + punto)
        NUM_PULSOS_TOP: positive := 5
    );

Port (     
           button_confir: in STD_LOGIC; --Confirmación de pedido
           vector_botones_monedas : in std_logic_vector (MONEDAS-1 downto 0);
           
           
           digsel : in STD_LOGIC_VECTOR (8 downto 0); --Los 9 productos que tenemos (switches)
           
           CLK    : in std_logic;
           RST    : in STD_LOGIC;
           digselec      : out std_logic_vector(NUM_DIGITS-1 downto 0);
           segment       : out STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
           
           ESTADO_OFF_button    : in STD_LOGIC;
           control_LEDS_1       : in STD_LOGIC;
           control_LEDS_2       : in STD_LOGIC;
           
           
           Err : out STD_LOGIC_VECTOR (15 downto 0)
           );
end TOP;

architecture Behavioral of TOP is
    
    signal clk_out : std_logic;
    
    -- SEÑALES DEL FSM
    signal estado_s       : unsigned(2 downto 0);
   
    
    -- SEÑALES MULTIPLEXOR     -------------------------------------------
    -- SEÑALES PARA LOS DIGITOS DEL DISPLAY, de tamaño 8 bits porque el último es el punto del dígito.
    -- Sirven como nexo entre el CTRL_DISPLAY y el Multiplexor que es quien se comunica con el HW
        signal DISP_DIG1_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG2_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG3_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG4_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG5_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG6_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG7_s    : std_logic_vector(NUM_SEGS-1 downto 0);
        signal DISP_DIG8_s    : std_logic_vector(NUM_SEGS-1 downto 0);  
    --Vector de los digitos síncrono, que permite al multiplexor decirle al HW qué digito activa por señal temporal
        signal dig_sel_sinc: STD_LOGIC_VECTOR (8 downto 0);
     
        
    -- Señales SINCRONIZADOR salida
    signal vector_productos_sinc       : std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
    signal vector_monedas_sinc         : std_logic_vector(Monedas-1 downto 0);
    signal boton_PAGO_sinc             : std_logic;

    -- Señales EDGEDTCTR salida
    signal edge_monedas_s              : std_logic;
    signal vector_monedas_deter_s      : std_logic_vector(Monedas-1 downto 0);
    signal edge_boton_pago_s           : std_logic;

    -- Señales Contador salida
    signal faltan_monedas_s : unsigned(3 downto 0);
    signal ok_s, error_s       : std_logic;    
        
    -- Señales STOCK salida
    signal productoOk_s     : std_logic;
    signal errorProducto_s  : std_logic;
    signal producto_id_s    : unsigned(3 downto 0);
    
    signal STOCK_producto_i_s :  std_logic_vector(NUM_PRODUCTOS-1 downto 0);
  
    signal en_leds : std_logic; ------------    ---------------------------------------------------------------------------------- OJO
    -- Señales Máquina de estados salida
    signal reset_general  : std_logic;


COMPONENT Prescaler
port(
        clk_in  : in  std_logic;   -- 100 MHz
        rst     : in  std_logic;   -- Reset síncrono
        clk_out : out std_logic    -- 16 kHz
    );
END COMPONENT;

COMPONENT Sincronizador
 Generic(
        NUM_PRODUCTOS: POSITIVE;
        NUM_MONEDAS: POSITIVE      
    );
 port(
        CLK: in std_logic;
        
        AS_PRODUCTOS: in std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
        AS_MONEDAS: in std_logic_vector (NUM_MONEDAS - 1 downto 0); 
        AS_CONFI : in std_logic;
               
        S_PRODUCTOS: out std_logic_vector (NUM_PRODUCTOS - 1 downto 0);
        S_MONEDAS: out std_logic_vector (NUM_MONEDAS - 1 downto 0);
        S_CONFI : out std_logic
    ); 
END COMPONENT;

component EDGEDTCTR is
        Generic(
            NUM_MONEDAS  : positive; 
            NUM_PULSOS   : positive 
        );
        Port(
            CLK : in STD_LOGIC;

            SYNC_IN_MONEDAS        : in STD_LOGIC_VECTOR (NUM_MONEDAS -1 downto 0);
            SYNC_IN_CONFIRMACION   : in STD_LOGIC;
            RESET_EDGE_DTC         : in STD_LOGIC;

            EDGE_MONEDAS_DETECTADO : out STD_LOGIC;
            EDGE_BOTON_PAGO        : out STD_LOGIC;

            Vector_monedas_deter   : out STD_LOGIC_VECTOR (NUM_MONEDAS -1 downto 0)
        );
    end component;

    component contador_monedas is
        port(
            clk            : in  std_logic;
            edge_monedas   : in  std_logic;
            edge_confir    : in  std_logic;
            monedas        : in  std_logic_vector(3 downto 0);
            estado         : in  unsigned(2 downto 0);
            Reset_Contador : in std_logic ;

            faltan_monedas_contador : out unsigned(3 downto 0);
            ok             : out std_logic;
            error          : out std_logic
        );
    end component;

component stock is
        generic (
            NUM_PRODUCTOS : positive := 9;
            PROD_BITS     : positive := 4
        );
        port(
            clk            : in  std_logic;
            estado         : in  unsigned(2 downto 0);
            productos      : in  std_logic_vector(NUM_PRODUCTOS-1 downto 0);
            error_pago     : in  std_logic;
            RESET_STOCK    : in  std_logic;
            Boton_Confirmar : in  std_logic;


            productoOk     : out std_logic;
            errorProducto  : out std_logic;
            producto_id    : out unsigned(PROD_BITS-1 downto 0);
            STOCK_producto_i   : out std_logic_vector(NUM_PRODUCTOS-1 downto 0)
  
        );
    end component;

COMPONENT Maq_Estados is
    Port(
            Error_producto      : in std_logic;
            Error_Pago          : in std_logic;
            OK_Pago             : in std_logic;
            OK_Producto         : in std_logic;
            RESET               : in std_logic;
            CLK                 : in std_logic;
            ESTADO_OFF          : in std_logic;
            
            RESET_SALIDA :  out std_logic;
            ESTADO_SALIDA : out unsigned(2 downto 0);
            LEDS : out STD_LOGIC_VECTOR (6 downto 0)

            );
END COMPONENT;

 component Multiplex is
        generic (
            NUM_DIGITS :positive ;
            NUM_SEGS   :positive 
        );
        port (
            clk           : in  STD_LOGIC;

            DISP_DIG1     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG2     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG3     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG4     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG5     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG6     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG7     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            DISP_DIG8     : in  STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);

            segment_mult  : out STD_LOGIC_VECTOR(NUM_SEGS-1 downto 0);
            digselec_mult : out STD_LOGIC_VECTOR(NUM_DIGITS-1 downto 0)
        );
end component;

 component ctr_display is
        generic(
            NUM_SEGS : positive
        );
        port(
            clk : in  std_logic;
            estado         : in  unsigned(2 downto 0);
            productos      : in  std_logic_vector(8 downto 0);
            faltan_monedas_ctrl_display : in  unsigned(3 downto 0);

            DISP_DIG1      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG2      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG3      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG4      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG5      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG6      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG7      : out std_logic_vector(NUM_SEGS-1 downto 0);
            DISP_DIG8      : out std_logic_vector(NUM_SEGS-1 downto 0)
        );
    end component;

    

    
begin

Inst_Prescaler : Prescaler
    port map(
        clk_in  => clk,
        rst    => rst,
        clk_out => clk_out
    );

   -- SINCRONIZADOR
	
Inst_Sincronizador : Sincronizador
        generic map(
            NUM_PRODUCTOS => NUM_PRODUCTOS,
            NUM_MONEDAS   => Monedas
        )
        port map(
            CLK          => clk_out,
            AS_PRODUCTOS => digsel,
            AS_MONEDAS   => vector_botones_monedas,
            AS_CONFI     => button_confir,
            S_PRODUCTOS  => dig_sel_sinc,
            S_MONEDAS    => vector_monedas_sinc,
            S_CONFI      => boton_PAGO_sinc
        );
        
    Inst_Maq_Estados : Maq_Estados
    Port Map(
            Error_producto  => errorProducto_s,
            Error_Pago      => error_s,
            OK_Pago         => ok_s,
            OK_Producto     => productoOk_s,
            RESET           => rst,
            CLK             => clk_out,
            ESTADO_OFF      => ESTADO_OFF_button,
            
            RESET_SALIDA    => reset_general,
            ESTADO_SALIDA   => estado_s,
            LEDS(0)         => Err(9),
            LEDS(1)         => Err(10),
            LEDS(2)         => Err(11),
            LEDS(3)         => Err(12),
            LEDS(4)         => Err(13),
            LEDS(5)         => Err(14),
            LEDS(6)         => Err(15)
            );
            
    -- EDGE DETECTOR
    inst_EDGE_DETECT : EDGEDTCTR
        generic map(
            NUM_MONEDAS => 4,
            NUM_PULSOS => NUM_PULSOS_TOP
        )
        port map(
            CLK                    => clk_out,           
            SYNC_IN_MONEDAS        => vector_monedas_sinc,
            SYNC_IN_CONFIRMACION   => boton_PAGO_sinc,
            RESET_EDGE_DTC         => reset_general,

            EDGE_MONEDAS_DETECTADO => edge_monedas_s,
            EDGE_BOTON_PAGO        => edge_boton_pago_s,
            Vector_monedas_deter   => vector_monedas_deter_s
        );

    -- CONTADOR MONEDAS
    Inst_Contador : contador_monedas
        port map(
            clk            => clk_out,
            edge_monedas   => edge_monedas_s,
            edge_confir    => edge_boton_pago_s,
            monedas        => vector_monedas_deter_s,
            estado         => estado_s,
            Reset_Contador => reset_general,
            
            faltan_monedas_contador => faltan_monedas_s,
            ok             => ok_s,
            error          => error_s
        );

        Inst_Stock : stock
        generic map(
            NUM_PRODUCTOS => 9,
            PROD_BITS     => 4
        )
        port map(
            clk            => clk_out,
            estado         => estado_s,
            productos      => dig_sel_sinc,
            error_pago     => error_s,
            RESET_STOCK    => reset_general,
            Boton_Confirmar => edge_boton_pago_s,


            productoOk     => productoOk_s,
            errorProducto  => errorProducto_s,
            producto_id    => producto_id_s,
            STOCK_producto_i => STOCK_producto_i_s
        );

    
    
    Inst_CTR_Display : ctr_display
        generic map(
            NUM_SEGS => NUM_SEGS
        )
        port map(
            clk            => clk_out,
            estado          => estado_s,
            productos       => dig_sel_sinc,
            faltan_monedas_ctrl_display  => faltan_monedas_s,

            DISP_DIG1       => DISP_DIG1_s,
            DISP_DIG2       => DISP_DIG2_s,
            DISP_DIG3       => DISP_DIG3_s,
            DISP_DIG4       => DISP_DIG4_s,
            DISP_DIG5       => DISP_DIG5_s,
            DISP_DIG6       => DISP_DIG6_s,
            DISP_DIG7       => DISP_DIG7_s,
            DISP_DIG8       => DISP_DIG8_s
        );
        
        
Inst_Multi : Multiplex
        generic map(
            NUM_DIGITS => NUM_DIGITS,
            NUM_SEGS   => NUM_SEGS
        )
        port map(
            clk           => clk_out,

            DISP_DIG1     => DISP_DIG1_s,
            DISP_DIG2     => DISP_DIG2_s,
            DISP_DIG3     => DISP_DIG3_s,
            DISP_DIG4     => DISP_DIG4_s,
            DISP_DIG5     => DISP_DIG5_s,
            DISP_DIG6     => DISP_DIG6_s,
            DISP_DIG7     => DISP_DIG7_s,
            DISP_DIG8     => DISP_DIG8_s,

            segment_mult  => segment,
            digselec_mult => digselec
        );
    



---Err(0) <= '1' when (estado_s /= 0) else '0';
--Err(1)  <=  dig_sel_sinc (0);
--Err(2)  <=  dig_sel_sinc (1);
--Err(3) <= error_s;

--Err(4) <= reset_general;
 
--Err(5)<= productoOk_s;
--Err(6)<= errorProducto_s;
--Err(7) <= '1' when (producto_id_s /= 0) else '0';

--PRUEBAS GUILLE

---- IF CONTROL DE LOS LEDS 1
--Err(0) <= STOCK_producto_i_s(0) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(1) <= STOCK_producto_i_s(1) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(2) <= STOCK_producto_i_s(2) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(3) <= STOCK_producto_i_s(3) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(4) <= STOCK_producto_i_s(4) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(5) <= STOCK_producto_i_s(5) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(6) <= STOCK_producto_i_s(6) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(7) <= STOCK_producto_i_s(7) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';
--Err(8) <= STOCK_producto_i_s(8) when (control_LEDS_1 = '1' and control_LEDS_2 = '0' ) else '0';


---- if  CONTROL DE LOS LEDS 2
--Err(0) <= STOCK_producto_i_s(0) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(1) <= STOCK_producto_i_s(1) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(2) <= STOCK_producto_i_s(2) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(3) <= STOCK_producto_i_s(3) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(4) <= STOCK_producto_i_s(4) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(5) <= STOCK_producto_i_s(5) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(6) <= STOCK_producto_i_s(6) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(7) <= STOCK_producto_i_s(7) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';
--Err(8) <= STOCK_producto_i_s(8) when (control_LEDS_2 = '1' and control_LEDS_1 = '0' ) else '0';


en_leds <= control_LEDS_1 xor control_LEDS_2;

Err(0) <= STOCK_producto_i_s(0) when en_leds = '1' else '0';
Err(1) <= STOCK_producto_i_s(1) when en_leds = '1' else '0';
Err(2) <= STOCK_producto_i_s(2) when en_leds = '1' else '0';
Err(3) <= STOCK_producto_i_s(3) when en_leds = '1' else '0';
Err(4) <= STOCK_producto_i_s(4) when en_leds = '1' else '0';
Err(5) <= STOCK_producto_i_s(5) when en_leds = '1' else '0';
Err(6) <= STOCK_producto_i_s(6) when en_leds = '1' else '0';
Err(7) <= STOCK_producto_i_s(7) when en_leds = '1' else '0';
Err(8) <= STOCK_producto_i_s(8) when en_leds = '1' else '0';

--Usaremos del Led 9 al 15 para mostrar que se está expendiendo 

-- MAS PRUEBAS
--Err(10) <= '1' when (errorProducto_s/= '0') else '0';  -- std_logig BIT


--Err(15) <= '1' when (estado_s = to_unsigned(0, estado_s'length)) else '0';
--Err(14) <= '1' when (estado_s = to_unsigned(1, estado_s'length)) else '0';
--Err(13) <= '1' when (estado_s = to_unsigned(2, estado_s'length)) else '0';
--Err(12) <= '1' when (estado_s = to_unsigned(3, estado_s'length)) else '0';
--Err(11) <= '1' when (estado_s = to_unsigned(4, estado_s'length)) else '0';

end Behavioral;


